-------------------------------------------------------------------
-- Name        : testbench.vhd
-- Author      : Enzzo Comassetto dos Santos
-- Version     : 0.1
-- Copyright   : Enzzo, Departamento de Eletrônica, Florianópolis, IFSC
-- Description : Script Modelsim para verificar o funcionamento do Contador de programa
-------------------------------------------------------------------

-- Bibliotecas e clásulas
LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
----------------------------------------------
ENTITY testbench IS
END ENTITY testbench;

ARCHITECTURE stimulus OF testbench IS
    -- Declaração de sinais
    signal clk        : std_logic; --Clock
    signal reset     : std_logic; --reset assícrono
    signal load    : std_logic; --Controle de escrita síncrono
    signal up       : std_logic; --Incrementa o valor do registrador
    signal datain     : std_logic_vector(15 downto 0); --Entrada de 16bits
    signal data    : std_logic_vector(15 downto 0); --Saida d 16 bits

BEGIN
    -- Instância do registrador
    dut : entity work.pc
        port map(
            clk     => clk,
            reset  => reset,
            load => load,
            up => up,
            datain  => datain,
            data => data
	
        );
    --Sequência de processos para verificar o funcionamento.
    process
    begin
        clk <= '0';
        wait for 10 ns;
        clk <= '1';
        wait for 10 ns;
    end process;

    Test : process
    begin
        reset  <= '1';
        load <= '0';
        up <= '0';
        datain  <= x"FFFF";
        wait for 60 ns;

        reset  <= '0';
        load <= '1';
        up <= '0';
        datain  <= x"FFFE";
        wait for 60 ns;

        reset  <= '0';
        load <= '1';
        up <= '1';
        datain  <= x"FFFD";
        wait for 60 ns;

        reset  <= '0';
        load <= '0';
        up <= '1';
        datain  <= x"FFFC";
        wait for 60 ns;

    end process Test;

END ARCHITECTURE stimulus;
